library ieee;
use ieee.std_logic_1164.all;
use work.pongtypes.all;

entity entity_number is
    port
    (
        number_pos_x_in     : in integer range 0 to 640;
        number_pos_y_in     : in integer range 0 to 480;

        number_start_x_in   : in integer range 0 to 640;
        number_start_y_in   : in integer range 0 to 480;
	
        number_score_in     : in score;


        number_colour_out   : out color
        );
end entity;


architecture architecture_number of entity_number is
    constant zero : number := ( ('0', '0', '1', '1', '1', '1', '0', '0'),
                                ('0', '1', '1', '0', '0', '1', '1', '0'),
                                ('1', '1', '0', '0', '0', '0', '1', '1'),
                                ('1', '1', '0', '0', '0', '0', '1', '1'),
                                ('1', '1', '0', '0', '0', '0', '1', '1'),
                                ('1', '1', '0', '0', '0', '0', '1', '1'),
                                ('1', '1', '0', '0', '0', '0', '1', '1'),
                                ('1', '1', '0', '0', '0', '0', '1', '1'),
                                ('1', '1', '0', '0', '0', '0', '1', '1'),
                                ('1', '1', '0', '0', '0', '0', '1', '1'),
                                ('0', '1', '1', '0', '0', '1', '1', '0'),
                                ('0', '0', '1', '1', '1', '1', '0', '0'));

    constant one : number := (  ('0', '0', '1', '1', '1', '0', '0', '0'),
                                ('1', '1', '1', '1', '1', '0', '0', '0'),
                                ('0', '0', '0', '1', '1', '0', '0', '0'),
                                ('0', '0', '0', '1', '1', '0', '0', '0'),
                                ('0', '0', '0', '1', '1', '0', '0', '0'),
                                ('0', '0', '0', '1', '1', '0', '0', '0'),
                                ('0', '0', '0', '1', '1', '0', '0', '0'),
                                ('0', '0', '0', '1', '1', '0', '0', '0'),
                                ('0', '0', '0', '1', '1', '0', '0', '0'),
                                ('0', '0', '0', '1', '1', '0', '0', '0'),
                                ('0', '0', '0', '1', '1', '0', '0', '0'),
                                ('1', '1', '1', '1', '1', '1', '1', '1'));

    constant two : number := (  ('0', '0', '1', '1', '1', '1', '0', '0'),
                                ('0', '1', '1', '0', '0', '1', '1', '0'),
                                ('1', '1', '0', '0', '0', '0', '1', '1'),
                                ('0', '0', '0', '0', '0', '0', '1', '1'),
                                ('0', '0', '0', '0', '0', '0', '1', '1'),
                                ('0', '0', '0', '0', '0', '1', '1', '0'),
                                ('0', '0', '0', '0', '1', '1', '0', '0'),
                                ('0', '0', '0', '1', '1', '0', '0', '0'),
                                ('0', '0', '1', '1', '0', '0', '0', '0'),
                                ('0', '1', '1', '0', '0', '0', '1', '1'),
                                ('1', '1', '0', '0', '0', '0', '1', '1'),
                                ('1', '1', '1', '1', '1', '1', '1', '1'));

    constant three : number := (('0', '1', '1', '1', '1', '1', '0', '0'),
                                ('1', '1', '0', '0', '0', '1', '1', '0'),
                                ('0', '0', '0', '0', '0', '0', '1', '1'),
                                ('0', '0', '0', '0', '0', '0', '1', '1'),
                                ('0', '0', '0', '0', '0', '1', '1', '0'),
                                ('0', '0', '0', '1', '1', '1', '0', '0'),
                                ('0', '0', '0', '0', '0', '1', '1', '0'),
                                ('0', '0', '0', '0', '0', '0', '1', '1'),
                                ('0', '0', '0', '0', '0', '0', '1', '1'),
                                ('0', '0', '0', '0', '0', '0', '1', '1'),
                                ('1', '1', '0', '0', '0', '1', '1', '0'),
                                ('0', '1', '1', '1', '1', '1', '0', '0'));

    constant four : number := ( ('0', '0', '0', '0', '0', '1', '1', '0'),
                                ('0', '0', '0', '0', '1', '1', '1', '0'),
                                ('0', '0', '0', '0', '1', '1', '1', '0'),
                                ('0', '0', '0', '1', '1', '1', '1', '0'),
                                ('0', '0', '1', '1', '0', '1', '1', '0'),
                                ('0', '0', '1', '1', '0', '1', '1', '0'),
                                ('0', '1', '1', '0', '0', '1', '1', '0'),
                                ('1', '1', '0', '0', '0', '1', '1', '0'),
                                ('1', '1', '1', '1', '1', '1', '1', '1'),
                                ('0', '0', '0', '0', '0', '1', '1', '0'),
                                ('0', '0', '0', '0', '0', '1', '1', '0'),
                                ('0', '0', '0', '1', '1', '1', '1', '1'));

    constant five : number := ( ('1', '1', '1', '1', '1', '1', '1', '0'),
                                ('1', '1', '0', '0', '0', '0', '0', '0'),
                                ('1', '1', '0', '0', '0', '0', '0', '0'),
                                ('1', '1', '0', '0', '0', '0', '0', '0'),
                                ('1', '1', '1', '1', '1', '1', '0', '0'),
                                ('1', '1', '0', '0', '0', '1', '1', '0'),
                                ('0', '0', '0', '0', '0', '0', '1', '1'),
                                ('0', '0', '0', '0', '0', '0', '1', '1'),
                                ('0', '0', '0', '0', '0', '0', '1', '1'),
                                ('0', '0', '0', '0', '0', '0', '1', '1'),
                                ('1', '1', '0', '0', '0', '1', '1', '0'),
                                ('0', '1', '1', '1', '1', '1', '0', '0'));

    constant six : number := (  ('0', '0', '0', '0', '1', '1', '1', '1'),
                                ('0', '0', '1', '1', '1', '0', '0', '0'),
                                ('0', '1', '1', '0', '0', '0', '0', '0'),
                                ('0', '1', '1', '0', '0', '0', '0', '0'),
                                ('1', '1', '0', '0', '0', '0', '0', '0'),
                                ('1', '1', '1', '1', '1', '1', '0', '0'),
                                ('1', '1', '1', '0', '0', '1', '1', '0'),
                                ('1', '1', '0', '0', '0', '0', '1', '1'),
                                ('1', '1', '0', '0', '0', '0', '1', '1'),
                                ('1', '1', '0', '0', '0', '0', '1', '1'),
                                ('0', '1', '1', '0', '0', '1', '1', '0'),
                                ('0', '0', '1', '1', '1', '1', '0', '0'));

    constant seven : number := (('1', '1', '1', '1', '1', '1', '1', '1'),
                                ('1', '1', '0', '0', '0', '0', '1', '1'),
                                ('1', '1', '0', '0', '0', '0', '1', '1'),
                                ('0', '0', '0', '0', '0', '1', '1', '0'),
                                ('0', '0', '0', '0', '0', '1', '1', '0'),
                                ('0', '0', '0', '0', '1', '1', '0', '0'),
                                ('0', '0', '0', '0', '1', '1', '0', '0'),
                                ('0', '0', '0', '1', '1', '0', '0', '0'),
                                ('0', '0', '0', '1', '1', '0', '0', '0'),
                                ('0', '0', '1', '1', '0', '0', '0', '0'),
                                ('0', '0', '1', '1', '0', '0', '0', '0'),
                                ('0', '0', '1', '1', '0', '0', '0', '0'));

    constant eight : number := (('0', '0', '1', '1', '1', '1', '0', '0'),
                                ('0', '1', '1', '0', '0', '1', '1', '0'),
                                ('1', '1', '0', '0', '0', '0', '1', '1'),
                                ('1', '1', '0', '0', '0', '0', '1', '1'),
                                ('0', '1', '1', '0', '0', '1', '1', '0'),
                                ('0', '0', '1', '1', '1', '1', '0', '0'),
                                ('0', '1', '1', '0', '0', '1', '1', '0'),
                                ('1', '1', '0', '0', '0', '0', '1', '1'),
                                ('1', '1', '0', '0', '0', '0', '1', '1'),
                                ('1', '1', '0', '0', '0', '0', '1', '1'),
                                ('0', '1', '1', '0', '0', '1', '1', '0'),
                                ('0', '0', '1', '1', '1', '1', '0', '0'));

    constant nine : number := ( ('0', '0', '1', '1', '1', '1', '0', '0'),
                                ('0', '1', '1', '0', '0', '1', '1', '0'),
                                ('1', '1', '0', '0', '0', '0', '1', '1'),
                                ('1', '1', '0', '0', '0', '0', '1', '1'),
                                ('1', '1', '0', '0', '0', '0', '1', '1'),
                                ('0', '1', '1', '0', '0', '1', '1', '1'),
                                ('0', '0', '1', '1', '1', '1', '1', '1'),
                                ('0', '0', '0', '0', '0', '0', '1', '1'),
                                ('0', '0', '0', '0', '0', '1', '1', '0'),
                                ('0', '0', '0', '0', '0', '1', '1', '0'),
                                ('0', '0', '0', '1', '1', '1', '0', '0'),
                                ('1', '1', '1', '1', '0', '0', '0', '0'));

    constant colour_max : color := (red => "1111", green => "1111", blue => "1111");
    constant colour_min : color := ("0000", "0000", "0000");
begin

    number_p : process(number_pos_x_in, number_pos_y_in)
    variable value      : integer range 0 to 9;
    variable num        : number;
    variable shift_x    : integer range 0 to 50 := 0;
    begin
        if(number_pos_x_in = 0 or number_pos_y_in = 0) then
            number_colour_out <= colour_min;
        else

        	shift_x := 0;

		    for i in 0 to 3 loop
		        value := number_score_in(i);


		        if(value = 0) then
		            num := zero;
		        elsif(value = 1) then
		            num := one;
		        elsif(value = 2) then
		            num := two;
		        elsif(value = 3) then
		            num := three;
		        elsif(value = 4) then
		            num := four;
		        elsif(value = 5) then
		            num := five;
		        elsif(value = 6) then
		            num := six;
		        elsif(value = 7) then
		            num := seven;
		        elsif(value = 8) then
		            num := eight;
		        else
		            num := nine;
		        end if;

		        if(number_pos_x_in >= number_start_x_in + shift_x and number_pos_y_in >= number_start_y_in and number_pos_x_in < number_start_x_in + 8 + shift_x and number_pos_y_in < number_start_y_in + 12) then
		            if(num(number_pos_y_in - number_start_y_in, number_pos_x_in - number_start_x_in) = '1') then
		                number_colour_out <= colour_max;
		                exit;
		            else
		                number_colour_out <= colour_min;
		                exit;
		            end if;
		        else
		            number_colour_out <= colour_min;
		        end if;
	        end loop;
        end if;
    end process;
end architecture architecture_number;
