

entity entity_pixelgenerator is
end entity;
